module load_to_mem(
    input bit clk,
    input bit rst_n,
    output reg[10:0] addr,
    output reg[9:0] data_out,
    output bit write_enable,
    input bit do_load,
    output bit did_load
);
    typedef enum {IDLE, START, LOOP, STORE, INCREMENT_INDEX, END} state_type;
    
    state_type state;

    const bit signed [9:0] noteA[0:1023] = {200, 0, 0, 200, 0, 200, 0, 200, 0, 200, 200, 0, 200, 0, 200, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 200, 200, 200, 200, 200, 0, 0, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 0, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 0, 0, 0, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 200, 0, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 200, 0, 0, 0, 200, 0, 0, 200, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0};
    const bit signed [9:0] noteB[0:1023] = {0, 200, 0, 200, 0, 200, 0, 0, 200, 0, 200, 0, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 200, 200, 0, 200, 0, 0, 200, 0, 200, 200, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 200, 200, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 0, 200, 0, 0, 200, 0, 0, 0, 200, 0, 0, 200, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 0, 200, 0, 200, 200, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 0, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 0, 200, 200, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 200, 200, 200, 0, 200, 0, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 200, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 200, 0, 0, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 0, 0, 0, 200, 200, 200, 200, 200, 0, 200, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200};
    const bit signed [9:0] noteD[0:1023] = {200, 0, 200, 0, 200, 200, 0, 200, 0, 200, 0, 200, 200, 0, 200, 0, 200, 0, 200, 0, 0, 200, 0, 200, 0, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 0, 0, 0, 0, 200, 200, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 0, 200, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 200, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 0, 0, 0, 0, 200, 0, 200, 200, 200, 0, 0, 200, 0, 0, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 0, 0, 0, 200, 200, 0, 200, 200, 0, 200, 0, 0, 0, 200, 0, 0, 200, 0, 200, 200, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 200, 200, 0, 200, 0, 0, 0, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 0, 0, 0, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 0, 0, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200};
    const bit signed [9:0] noteE[0:1023] = {200, 200, 0, 200, 0, 200, 0, 200, 200, 0, 200, 0, 200, 0, 200, 0, 0, 200, 0, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200};
    const bit signed [9:0] noteE2[0:1023] = {0, 200, 0, 200, 0, 200, 0, 0, 200, 0, 200, 0, 200, 0, 0, 200, 0, 200, 0, 200, 0, 200, 200, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 200, 0, 200, 200, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 200, 0, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 0, 200, 0, 0, 0, 0, 200, 200, 0, 200, 200, 200, 200, 200, 200, 0, 200, 200, 200, 0, 0, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 0, 0, 0, 0, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 0, 0, 0, 200, 0, 200, 0, 0, 0, 200, 200, 200, 200, 200, 200, 0, 0, 200, 0, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 0, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 200, 200, 200, 200, 0, 0, 200, 0, 0, 0, 0, 200, 200, 0, 200, 200, 0, 200, 200, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 0, 0, 0, 200, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200};
    const bit signed [9:0] noteG[0:1023] = {200, 0, 0, 200, 0, 200, 0, 200, 0, 200, 200, 0, 200, 0, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 200, 200, 0, 200, 200, 200, 0, 0, 0, 0, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 200, 200, 200, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 0, 200, 200, 0, 0, 200, 200, 0, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 0, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 0, 200, 200, 200, 200, 0, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 200, 200, 200, 200, 200, 0, 0, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 0, 0, 200, 200, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 0, 0, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 0, 200, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 200, 200, 200, 200, 0, 0, 0, 0, 0, 0, 0, 200, 0, 200, 200, 200, 0, 200, 0, 0, 200, 0, 0, 200, 200, 0, 0, 200, 0, 0, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 0, 200, 0, 0, 200, 0, 200, 0, 0, 200, 200, 0, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 0, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 200, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 0, 0, 200, 200, 200, 200, 0, 200, 200, 200, 200, 0, 0, 200, 0, 200, 0, 0, 200, 200, 200, 0, 0, 200};
    const bit signed [9:0] noteE2_2[0:1023] = {4, 59, 30, 16, 20, 54, 4, 8, 61, 2, 4, 60, 59, 6, 57, 55, 3, 59, 53, 3, 1, 60, 6, 4, 60, 9, 5, 57, 63, 4, 58, 7, 11, 57, 63, 2, 53, 61, 61, 56, 60, 2, 1, 0, 8, 63, 63, 9, 62, 59, 7, 60, 57, 2, 59, 56, 0, 62, 57, 5, 6, 60, 4, 5, 60, 4, 5, 56, 0, 4, 58, 1, 2, 58, 0, 5, 63, 63, 7, 0, 1, 8, 62, 62, 8, 63, 63, 6, 0, 62, 7, 2, 55, 4, 3, 60, 9, 63, 53, 1, 58, 50, 58, 63, 57, 63, 4, 57, 62, 5, 61, 0, 4, 59, 2, 6, 62, 59, 2, 59, 56, 62, 62, 61, 9, 7, 56, 6, 2, 53, 4, 59, 52, 1, 63, 62, 4, 3, 61, 1, 8, 61, 61, 5, 53, 61, 3, 59, 4, 5, 63, 63, 2, 59, 56, 2, 59, 58, 6, 60, 59, 3, 60, 57, 3, 1, 59, 6, 4, 59, 5, 3, 57, 2, 3, 58, 1, 4, 58, 62, 2, 56, 61, 2, 60, 63, 4, 62, 63, 6, 61, 61, 6, 63, 61, 7, 63, 60, 4, 63, 57, 2, 0, 56, 2, 0, 56, 1, 2, 58, 2, 4, 60, 1, 5, 60, 63, 4, 59, 63, 3, 60, 61, 2, 59, 59, 3, 59, 60, 5, 63, 61, 6, 0, 62, 6, 3, 59, 5, 2, 57, 4, 1, 56, 1, 2, 58, 0, 3, 59, 63, 4, 59, 63, 4, 59, 63, 4, 61, 62, 4, 61, 61, 5, 60, 60, 4, 61, 58, 3, 63, 58, 3, 1, 57, 4, 3, 58, 3, 4, 58, 3, 4, 59, 1, 4, 59, 63, 4, 59, 62, 3, 59, 62, 4, 61, 62, 6, 62, 62, 6, 62, 60, 5, 63, 59, 3, 0, 58, 3, 1, 58, 2, 2, 57, 2, 3, 59, 1, 3, 59, 0, 4, 60, 63, 4, 59, 62, 3, 60, 62, 3, 62, 60, 5, 62, 60, 5, 62, 59, 4, 0, 59, 3, 2, 59, 2, 3, 58, 2, 3, 58, 0, 3, 58, 63, 4, 60, 63, 5, 61, 62, 4, 61, 61, 3, 63, 61, 4, 63, 60, 2, 63, 59, 2, 0, 59, 2, 1, 60, 1, 3, 59, 1, 4, 59, 1, 3, 59, 0, 4, 59, 63, 4, 61, 62, 3, 60, 62, 3, 61, 62, 3, 62, 62, 3, 63, 62, 4, 63, 60, 3, 0, 60, 3, 0, 60, 2, 2, 59, 1, 2, 59, 1, 3, 59, 1, 3, 60, 0, 4, 61, 63, 4, 61, 63, 3, 61, 62, 3, 61, 61, 3, 63, 61, 3, 63, 61, 3, 0, 60, 2, 1, 60, 2, 3, 59, 1, 3, 60, 1, 2, 59, 0, 3, 60, 63, 3, 61, 63, 4, 61, 62, 3, 62, 61, 3, 62, 61, 3, 62, 60, 3, 0, 59, 2, 0, 59, 2, 1, 59, 2, 2, 59, 1, 2, 59, 2, 3, 60, 0, 3, 60, 63, 3, 60, 62, 3, 61, 62, 3, 61, 62, 4, 62, 61, 3, 63, 60, 3, 63, 61, 3, 1, 59, 2, 3, 60, 2, 2, 59, 2, 3, 59, 0, 3, 60, 0, 3, 60, 63, 4, 60, 63, 3, 62, 62, 3, 61, 61, 3, 62, 61, 3, 63, 61, 3, 1, 60, 2, 2, 60, 2, 2, 59, 2, 3, 59, 0, 2, 60, 0, 3, 60, 0, 3, 60, 62, 2, 60, 62, 2, 61, 61, 2, 62, 61, 2, 63, 60, 2, 0, 60, 1, 0, 59, 1, 2, 58, 1, 3, 59, 1, 2, 59, 0, 3, 60, 63, 4, 61, 63, 3, 61, 62, 2, 62, 62, 2, 62, 61, 2, 63, 61, 2, 1, 60, 3, 1, 60, 2, 2, 59, 2, 2, 59, 2, 3, 60, 0, 2, 60, 63, 3, 60, 63, 3, 61, 62, 2, 61, 62, 3, 62, 61, 3, 62, 60, 2, 0, 60, 2, 0, 61, 2, 1, 60, 2, 3, 60, 1, 2, 60, 1, 3, 61, 1, 3, 61, 63, 2, 61, 63, 3, 62, 62, 3, 62, 61, 2, 62, 61, 2, 63, 61, 1, 0, 60, 2, 0, 60, 1, 1, 60, 0, 1, 60, 1, 2, 60, 0, 2, 60, 63, 1, 61, 62, 2, 62, 63, 2, 62, 62, 2, 63, 61, 1, 63, 62, 2, 0, 61, 2, 0, 61, 1, 1, 62, 1, 2, 61, 1, 2, 61, 0, 3, 61, 1, 2, 61, 63, 2, 61, 63, 2, 61, 63, 2, 62, 61, 2, 62, 62, 1, 63, 61, 2, 0, 61, 1, 0, 62, 1, 1, 61, 0, 2, 61, 0, 2, 61, 0, 2, 61, 0, 2, 62, 0, 2, 62, 63, 2, 62, 63, 2, 63, 63, 1, 63, 63, 1, 63, 62, 2, 63, 62, 1, 0, 61, 0, 1, 61, 0, 2, 61, 1, 2, 60, 63, 2, 61, 63, 2, 61, 63, 2, 61, 63, 2, 62, 63, 1, 62, 63, 1, 63, 63, 1, 0, 62, 1, 0, 62, 1, 1, 62, 1, 1, 61, 1, 2, 61, 1, 2, 61, 0, 2, 62, 0, 1, 62, 63, 1, 62, 63, 1, 62, 63, 1, 63, 62, 1, 0, 62, 1, 0, 61, 1, 0, 62, 0, 1, 61, 0, 1, 62, 0, 1, 62, 0, 1, 62, 0, 2, 62, 0, 0, 62, 0, 2, 63, 63, 1, 62, 63, 1, 63, 63, 1, 0, 62, 0, 0, 62, 1, 0, 62, 0, 0, 61, 0, 1, 61, 0, 1, 61, 63, 1, 61, 0, 0, 62, 63, 1, 63, 63, 1, 62, 63, 1, 62, 63, 1, 63, 63, 2, 63, 63, 1, 0, 62, 1, 0, 62, 0, 1, 62, 0, 2, 62, 0, 1, 62, 0, 1, 62, 63, 1, 62, 63, 1, 62, 63, 1, 63, 63, 1, 63, 63, 1, 63, 62, 0, 0, 63, 0, 63, 62, 1, 0, 62, 0, 0, 62, 0, 0, 62, 0, 1, 62, 0, 1, 62, 0, 1, 63, 0, 1, 63, 0, 1, 63, 63, 1, 63, 63, 1, 63, 63, 1, 63, 62, 1, 0};
    
    reg [10:0] index;
    wire [10:0] index_inv;
    assign index_inv[0] = index[9];
    assign index_inv[1] = index[8];
    assign index_inv[2] = index[7];
    assign index_inv[3] = index[6];
    assign index_inv[4] = index[5];
    assign index_inv[5] = index[4];
    assign index_inv[6] = index[3];
    assign index_inv[7] = index[2];
    assign index_inv[8] = index[1];
    assign index_inv[9] = index[0];
    assign index_inv[10] = 0;

    always @(posedge clk) begin
        if(rst_n == 0) begin
            state <= IDLE;
            did_load <= 0;
        end else begin
            case(state)
                IDLE: begin
                    state <= START;
                end
                START: begin
                    index <= 0;
                    if(do_load == 1) begin
                        state <= LOOP;                        
                    end else begin
                        state <= START;
                    end
                end
                LOOP: begin
                    if(index < 1024) begin
                        state <= STORE;
                    end else begin
                        state <= END;
                    end
                end
                STORE: begin
                    data_out <= noteE2_2[index];
                    addr <= index_inv;
                    write_enable <= 1;
                    state <= INCREMENT_INDEX;
                end
                INCREMENT_INDEX: begin
                    write_enable <= 0;
                    index <= index + 1;
                    state <= LOOP;
                end
                END: begin
                    state <= END;
                    did_load <= 1;
                end
            endcase
        end
    end


endmodule