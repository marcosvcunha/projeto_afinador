
module fft #(
        parameter N_bits=16, // N�mero de bits utilizados
        parameter SAMPLE_SIZE=1024 // Tamanho do 
)(
    input bit clk,
    input bit rst_n,
    output reg [10:0] addr,
    output bit write_enable,
    input wire [9:0] data_in,
    output wire [9:0] data_out_wire,
    input bit do_fft,
    output bit fft_done
);
    typedef enum {IDLE, START, LOOP_1, LOOP_2, LOOP_3, SET_ADDR, WAIT_DATA1, READ_MEM1, WAIT_DATA2, 
        READ_MEM2, WAIT_DATA3, READ_MEM3, WAIT_DATA4, READ_MEM4, MULT1, MULT2, MULT3, MULT4, DIV, 
        STORE1, STORE2, STORE3, STORE4, END} state_type;
    
    const bit signed [9:0] WnR[0:1023] = {511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 510, 510, 510, 510, 509, 509, 509, 508, 508, 508, 507, 507, 506, 506, 505, 505, 504, 504, 503, 503, 502, 502, 501, 500, 500, 499, 498, 498, 497, 496, 495, 495, 494, 493, 492, 491, 490, 489, 489, 488, 487, 486, 485, 484, 483, 482, 481, 479, 478, 477, 476, 475, 474, 473, 471, 470, 469, 468, 466, 465, 464, 462, 461, 460, 458, 457, 455, 454, 453, 451, 450, 448, 447, 445, 443, 442, 440, 439, 437, 435, 434, 432, 430, 429, 427, 425, 423, 422, 420, 418, 416, 414, 413, 411, 409, 407, 405, 403, 401, 399, 397, 395, 393, 391, 389, 387, 385, 383, 381, 379, 377, 375, 372, 370, 368, 366, 364, 362, 359, 357, 355, 353, 350, 348, 346, 343, 341, 339, 336, 334, 332, 329, 327, 324, 322, 319, 317, 314, 312, 310, 307, 304, 302, 299, 297, 294, 292, 289, 287, 284, 281, 279, 276, 273, 271, 268, 265, 263, 260, 257, 255, 252, 249, 246, 244, 241, 238, 235, 233, 230, 227, 224, 221, 218, 216, 213, 210, 207, 204, 201, 198, 195, 193, 190, 187, 184, 181, 178, 175, 172, 169, 166, 163, 160, 157, 154, 151, 148, 145, 142, 139, 136, 133, 130, 127, 124, 121, 118, 115, 112, 109, 106, 102, 99, 96, 93, 90, 87, 84, 81, 78, 75, 72, 68, 65, 62, 59, 56, 53, 50, 47, 43, 40, 37, 34, 31, 28, 25, 21, 18, 15, 12, 9, 6, 3, 0, -3, -6, -9, -12, -15, -18, -21, -25, -28, -31, -34, -37, -40, -43, -47, -50, -53, -56, -59, -62, -65, -68, -72, -75, -78, -81, -84, -87, -90, -93, -96, -99, -102, -106, -109, -112, -115, -118, -121, -124, -127, -130, -133, -136, -139, -142, -145, -148, -151, -154, -157, -160, -163, -166, -169, -172, -175, -178, -181, -184, -187, -190, -193, -195, -198, -201, -204, -207, -210, -213, -216, -218, -221, -224, -227, -230, -233, -235, -238, -241, -244, -246, -249, -252, -255, -257, -260, -263, -265, -268, -271, -273, -276, -279, -281, -284, -287, -289, -292, -294, -297, -299, -302, -304, -307, -310, -312, -314, -317, -319, -322, -324, -327, -329, -332, -334, -336, -339, -341, -343, -346, -348, -350, -353, -355, -357, -359, -362, -364, -366, -368, -370, -372, -375, -377, -379, -381, -383, -385, -387, -389, -391, -393, -395, -397, -399, -401, -403, -405, -407, -409, -411, -413, -414, -416, -418, -420, -422, -423, -425, -427, -429, -430, -432, -434, -435, -437, -439, -440, -442, -443, -445, -447, -448, -450, -451, -453, -454, -455, -457, -458, -460, -461, -462, -464, -465, -466, -468, -469, -470, -471, -473, -474, -475, -476, -477, -478, -479, -481, -482, -483, -484, -485, -486, -487, -488, -489, -489, -490, -491, -492, -493, -494, -495, -495, -496, -497, -498, -498, -499, -500, -500, -501, -502, -502, -503, -503, -504, -504, -505, -505, -506, -506, -507, -507, -508, -508, -508, -509, -509, -509, -510, -510, -510, -510, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -510, -510, -510, -510, -509, -509, -509, -508, -508, -508, -507, -507, -506, -506, -505, -505, -504, -504, -503, -503, -502, -502, -501, -500, -500, -499, -498, -498, -497, -496, -495, -495, -494, -493, -492, -491, -490, -489, -489, -488, -487, -486, -485, -484, -483, -482, -481, -479, -478, -477, -476, -475, -474, -473, -471, -470, -469, -468, -466, -465, -464, -462, -461, -460, -458, -457, -455, -454, -453, -451, -450, -448, -447, -445, -443, -442, -440, -439, -437, -435, -434, -432, -430, -429, -427, -425, -423, -422, -420, -418, -416, -414, -413, -411, -409, -407, -405, -403, -401, -399, -397, -395, -393, -391, -389, -387, -385, -383, -381, -379, -377, -375, -372, -370, -368, -366, -364, -362, -359, -357, -355, -353, -350, -348, -346, -343, -341, -339, -336, -334, -332, -329, -327, -324, -322, -319, -317, -314, -312, -310, -307, -304, -302, -299, -297, -294, -292, -289, -287, -284, -281, -279, -276, -273, -271, -268, -265, -263, -260, -257, -255, -252, -249, -246, -244, -241, -238, -235, -233, -230, -227, -224, -221, -218, -216, -213, -210, -207, -204, -201, -198, -195, -193, -190, -187, -184, -181, -178, -175, -172, -169, -166, -163, -160, -157, -154, -151, -148, -145, -142, -139, -136, -133, -130, -127, -124, -121, -118, -115, -112, -109, -106, -102, -99, -96, -93, -90, -87, -84, -81, -78, -75, -72, -68, -65, -62, -59, -56, -53, -50, -47, -43, -40, -37, -34, -31, -28, -25, -21, -18, -15, -12, -9, -6, -3, 0, 3, 6, 9, 12, 15, 18, 21, 25, 28, 31, 34, 37, 40, 43, 47, 50, 53, 56, 59, 62, 65, 68, 72, 75, 78, 81, 84, 87, 90, 93, 96, 99, 102, 106, 109, 112, 115, 118, 121, 124, 127, 130, 133, 136, 139, 142, 145, 148, 151, 154, 157, 160, 163, 166, 169, 172, 175, 178, 181, 184, 187, 190, 193, 195, 198, 201, 204, 207, 210, 213, 216, 218, 221, 224, 227, 230, 233, 235, 238, 241, 244, 246, 249, 252, 255, 257, 260, 263, 265, 268, 271, 273, 276, 279, 281, 284, 287, 289, 292, 294, 297, 299, 302, 304, 307, 310, 312, 314, 317, 319, 322, 324, 327, 329, 332, 334, 336, 339, 341, 343, 346, 348, 350, 353, 355, 357, 359, 362, 364, 366, 368, 370, 372, 375, 377, 379, 381, 383, 385, 387, 389, 391, 393, 395, 397, 399, 401, 403, 405, 407, 409, 411, 413, 414, 416, 418, 420, 422, 423, 425, 427, 429, 430, 432, 434, 435, 437, 439, 440, 442, 443, 445, 447, 448, 450, 451, 453, 454, 455, 457, 458, 460, 461, 462, 464, 465, 466, 468, 469, 470, 471, 473, 474, 475, 476, 477, 478, 479, 481, 482, 483, 484, 485, 486, 487, 488, 489, 489, 490, 491, 492, 493, 494, 495, 495, 496, 497, 498, 498, 499, 500, 500, 501, 502, 502, 503, 503, 504, 504, 505, 505, 506, 506, 507, 507, 508, 508, 508, 509, 509, 509, 510, 510, 510, 510, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511};
    const bit signed [9:0] WnI[0:1023] = {0, 3, 6, 9, 12, 15, 18, 21, 25, 28, 31, 34, 37, 40, 43, 47, 50, 53, 56, 59, 62, 65, 68, 72, 75, 78, 81, 84, 87, 90, 93, 96, 99, 102, 106, 109, 112, 115, 118, 121, 124, 127, 130, 133, 136, 139, 142, 145, 148, 151, 154, 157, 160, 163, 166, 169, 172, 175, 178, 181, 184, 187, 190, 193, 195, 198, 201, 204, 207, 210, 213, 216, 218, 221, 224, 227, 230, 233, 235, 238, 241, 244, 246, 249, 252, 255, 257, 260, 263, 265, 268, 271, 273, 276, 279, 281, 284, 287, 289, 292, 294, 297, 299, 302, 304, 307, 310, 312, 314, 317, 319, 322, 324, 327, 329, 332, 334, 336, 339, 341, 343, 346, 348, 350, 353, 355, 357, 359, 362, 364, 366, 368, 370, 372, 375, 377, 379, 381, 383, 385, 387, 389, 391, 393, 395, 397, 399, 401, 403, 405, 407, 409, 411, 413, 414, 416, 418, 420, 422, 423, 425, 427, 429, 430, 432, 434, 435, 437, 439, 440, 442, 443, 445, 447, 448, 450, 451, 453, 454, 455, 457, 458, 460, 461, 462, 464, 465, 466, 468, 469, 470, 471, 473, 474, 475, 476, 477, 478, 479, 481, 482, 483, 484, 485, 486, 487, 488, 489, 489, 490, 491, 492, 493, 494, 495, 495, 496, 497, 498, 498, 499, 500, 500, 501, 502, 502, 503, 503, 504, 504, 505, 505, 506, 506, 507, 507, 508, 508, 508, 509, 509, 509, 510, 510, 510, 510, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 511, 510, 510, 510, 510, 509, 509, 509, 508, 508, 508, 507, 507, 506, 506, 505, 505, 504, 504, 503, 503, 502, 502, 501, 500, 500, 499, 498, 498, 497, 496, 495, 495, 494, 493, 492, 491, 490, 489, 489, 488, 487, 486, 485, 484, 483, 482, 481, 479, 478, 477, 476, 475, 474, 473, 471, 470, 469, 468, 466, 465, 464, 462, 461, 460, 458, 457, 455, 454, 453, 451, 450, 448, 447, 445, 443, 442, 440, 439, 437, 435, 434, 432, 430, 429, 427, 425, 423, 422, 420, 418, 416, 414, 413, 411, 409, 407, 405, 403, 401, 399, 397, 395, 393, 391, 389, 387, 385, 383, 381, 379, 377, 375, 372, 370, 368, 366, 364, 362, 359, 357, 355, 353, 350, 348, 346, 343, 341, 339, 336, 334, 332, 329, 327, 324, 322, 319, 317, 314, 312, 310, 307, 304, 302, 299, 297, 294, 292, 289, 287, 284, 281, 279, 276, 273, 271, 268, 265, 263, 260, 257, 255, 252, 249, 246, 244, 241, 238, 235, 233, 230, 227, 224, 221, 218, 216, 213, 210, 207, 204, 201, 198, 195, 193, 190, 187, 184, 181, 178, 175, 172, 169, 166, 163, 160, 157, 154, 151, 148, 145, 142, 139, 136, 133, 130, 127, 124, 121, 118, 115, 112, 109, 106, 102, 99, 96, 93, 90, 87, 84, 81, 78, 75, 72, 68, 65, 62, 59, 56, 53, 50, 47, 43, 40, 37, 34, 31, 28, 25, 21, 18, 15, 12, 9, 6, 3, 0, -3, -6, -9, -12, -15, -18, -21, -25, -28, -31, -34, -37, -40, -43, -47, -50, -53, -56, -59, -62, -65, -68, -72, -75, -78, -81, -84, -87, -90, -93, -96, -99, -102, -106, -109, -112, -115, -118, -121, -124, -127, -130, -133, -136, -139, -142, -145, -148, -151, -154, -157, -160, -163, -166, -169, -172, -175, -178, -181, -184, -187, -190, -193, -195, -198, -201, -204, -207, -210, -213, -216, -218, -221, -224, -227, -230, -233, -235, -238, -241, -244, -246, -249, -252, -255, -257, -260, -263, -265, -268, -271, -273, -276, -279, -281, -284, -287, -289, -292, -294, -297, -299, -302, -304, -307, -310, -312, -314, -317, -319, -322, -324, -327, -329, -332, -334, -336, -339, -341, -343, -346, -348, -350, -353, -355, -357, -359, -362, -364, -366, -368, -370, -372, -375, -377, -379, -381, -383, -385, -387, -389, -391, -393, -395, -397, -399, -401, -403, -405, -407, -409, -411, -413, -414, -416, -418, -420, -422, -423, -425, -427, -429, -430, -432, -434, -435, -437, -439, -440, -442, -443, -445, -447, -448, -450, -451, -453, -454, -455, -457, -458, -460, -461, -462, -464, -465, -466, -468, -469, -470, -471, -473, -474, -475, -476, -477, -478, -479, -481, -482, -483, -484, -485, -486, -487, -488, -489, -489, -490, -491, -492, -493, -494, -495, -495, -496, -497, -498, -498, -499, -500, -500, -501, -502, -502, -503, -503, -504, -504, -505, -505, -506, -506, -507, -507, -508, -508, -508, -509, -509, -509, -510, -510, -510, -510, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -511, -510, -510, -510, -510, -509, -509, -509, -508, -508, -508, -507, -507, -506, -506, -505, -505, -504, -504, -503, -503, -502, -502, -501, -500, -500, -499, -498, -498, -497, -496, -495, -495, -494, -493, -492, -491, -490, -489, -489, -488, -487, -486, -485, -484, -483, -482, -481, -479, -478, -477, -476, -475, -474, -473, -471, -470, -469, -468, -466, -465, -464, -462, -461, -460, -458, -457, -455, -454, -453, -451, -450, -448, -447, -445, -443, -442, -440, -439, -437, -435, -434, -432, -430, -429, -427, -425, -423, -422, -420, -418, -416, -414, -413, -411, -409, -407, -405, -403, -401, -399, -397, -395, -393, -391, -389, -387, -385, -383, -381, -379, -377, -375, -372, -370, -368, -366, -364, -362, -359, -357, -355, -353, -350, -348, -346, -343, -341, -339, -336, -334, -332, -329, -327, -324, -322, -319, -317, -314, -312, -310, -307, -304, -302, -299, -297, -294, -292, -289, -287, -284, -281, -279, -276, -273, -271, -268, -265, -263, -260, -257, -255, -252, -249, -246, -244, -241, -238, -235, -233, -230, -227, -224, -221, -218, -216, -213, -210, -207, -204, -201, -198, -195, -193, -190, -187, -184, -181, -178, -175, -172, -169, -166, -163, -160, -157, -154, -151, -148, -145, -142, -139, -136, -133, -130, -127, -124, -121, -118, -115, -112, -109, -106, -102, -99, -96, -93, -90, -87, -84, -81, -78, -75, -72, -68, -65, -62, -59, -56, -53, -50, -47, -43, -40, -37, -34, -31, -28, -25, -21, -18, -15, -12, -9, -6, -3};

    reg signed [9:0] WnR_op;
    reg signed [9:0] WnI_op;

    state_type state;
    reg [3:0] LOOP_1_Counter; // Conta os estágios. Para 1024 amostras, vai de 0 a 9.
    reg [9:0] Nb; // Número de borboletas do estágio.
    reg [9:0] Np; // Número de "asas" na borboleta.
    reg [9:0] idxB; // Index de "cima" da borboleta.
    reg [8:0] Diff; // Variação dos index dos Omegas.
    reg [9:0] LOOP_2_Counter; // Conta o index das borboletas. O limite altera conforme o estado. (p/ 1024 amostras o máximo é 512) 
    reg [9:0] idx; // Index da saída atual a ser calculada
    reg [9:0] Widx; // Idx do Omega a ser usado
    reg [9:0] LOOP_3_Counter; // Conta o index da "asa" borboletas. (p/ 1024 amostras o máximo é 512)
    reg [9:0] idxCima;
    // wire [9:0] idxCima_inv;
    reg [9:0] idxBaixo;
    // wire [9:0] idxBaixo_inv;
    reg [9:0] data_out;
    
    assign data_out_wire = data_out;

    // assign idxCima_inv[0] = idxCima[9];
    // assign idxCima_inv[1] = idxCima[8];
    // assign idxCima_inv[2] = idxCima[7];
    // assign idxCima_inv[3] = idxCima[6];
    // assign idxCima_inv[4] = idxCima[5];
    // assign idxCima_inv[5] = idxCima[4];
    // assign idxCima_inv[6] = idxCima[3];
    // assign idxCima_inv[7] = idxCima[2];
    // assign idxCima_inv[8] = idxCima[1];
    // assign idxCima_inv[9] = idxCima[0];

    // assign idxBaixo_inv[0] = idxBaixo[9];
    // assign idxBaixo_inv[1] = idxBaixo[8];
    // assign idxBaixo_inv[2] = idxBaixo[7];
    // assign idxBaixo_inv[3] = idxBaixo[6];
    // assign idxBaixo_inv[4] = idxBaixo[5];
    // assign idxBaixo_inv[5] = idxBaixo[4];
    // assign idxBaixo_inv[6] = idxBaixo[3];
    // assign idxBaixo_inv[7] = idxBaixo[2];
    // assign idxBaixo_inv[8] = idxBaixo[1];
    // assign idxBaixo_inv[9] = idxBaixo[0];

    
    reg signed [9:0] fftRC; // Número Real de Cima 
    reg signed [9:0] fftIC; // Número Imaginário de Cima
    reg signed [9:0] fftRB; // Número Real de Baixo
    reg signed [9:0] fftIB; // Número Imaginário de Baixo

    reg signed [9:0] tempR;
    reg signed [9:0] tempI;

    wire signed [9:0] temp2R;
    reg signed [18:0] temp2R_aux;
    wire signed [9:0] temp2I;
    reg signed [18:0] temp2I_aux;
    int debug_count = 0;
    
    assign temp2R = temp2R_aux[18:9];
    assign temp2I = temp2I_aux[18:9];


    function reg[8:0] calc_diff(input reg [3:0] stage);
        case(stage)
            4'd0:
                calc_diff = 9'd0;
            4'd1:
                calc_diff = 9'd256;
            4'd2:
                calc_diff = 9'd128;
            4'd3:
                calc_diff = 9'd64;
            4'd4:
                calc_diff = 9'd32;
            4'd5:
                calc_diff = 9'd16;
            4'd6:
                calc_diff = 9'd8;
            4'd7:
                calc_diff = 9'd4;
            4'd8:
                calc_diff = 9'd2;
            4'd9:
                calc_diff = 9'd1;
        endcase
    endfunction



    always @(posedge clk) begin
        if(rst_n == 0 || do_fft == 0) begin
            state <= IDLE;
            fft_done <= 0;
            write_enable <= 0;
        end else begin
            case(state)
                IDLE:
                    begin
                        state <= START;
                        write_enable <= 0;
                    end
                START: begin
                    // TODO: puxar a entrada para a parte da memória relativa a parte real da transformada
                    LOOP_1_Counter <= 10'd0;
                    state <= LOOP_1;
                end
                LOOP_1:
                    if(LOOP_1_Counter == 4'd10) begin
                        state <= END;
                    end else begin
                        if(LOOP_1_Counter == 4'b0) begin
                            Nb <= 10'd512;
                            Np <= 10'd1;
                        end else begin
                            Nb <= Nb >> 1;
                            Np <= Np << 1;
                        end
                        Diff <= calc_diff(LOOP_1_Counter);
                        idxB <= 10'd0;
                        LOOP_1_Counter <= LOOP_1_Counter + 1;
                        LOOP_2_Counter <= 0;
                        state <= LOOP_2;
                    end
                LOOP_2:
                    if(LOOP_2_Counter == Nb) begin
                        state <= LOOP_1;
                    end else begin
                        idx <= idxB;
                        idxB <= idxB + (Np << 1);
                        Widx <= 10'd0;
                        LOOP_2_Counter <= LOOP_2_Counter + 1;
                        LOOP_3_Counter <= 0;
                        state <= LOOP_3;
                    end
                LOOP_3:
                    begin
                        write_enable <= 0;
                        if(LOOP_3_Counter == Np) begin
                            state <= LOOP_2;
                        end else begin
                            // Seta os endereços
                            idxCima <= idx;
                            idxBaixo <= idx + Np;
                            WnR_op <= WnR[Widx];
                            WnI_op <= WnI[Widx];
                            Widx <= Widx + Diff;
                            idx <= idx + 1;
                            LOOP_3_Counter <= LOOP_3_Counter + 1;
                            state <= SET_ADDR;
                        end
                    end
                SET_ADDR:
                    begin
                        addr <= idxCima;
                        state <= WAIT_DATA1;
                    end
                WAIT_DATA1:
                    state <= READ_MEM1;
                READ_MEM1:
                    begin
                        fftRC <= data_in;
                        tempR <= data_in;
                        addr <= idxCima + 1024;
                        state <= WAIT_DATA2;
                    end
                WAIT_DATA2:
                    state <= READ_MEM2;
                READ_MEM2:
                    begin
                        fftIC <= data_in;
                        tempI <= data_in;
                        addr <= idxBaixo;
                        state <= WAIT_DATA3;
                    end
                WAIT_DATA3:
                    state <= READ_MEM3;
                READ_MEM3:
                    begin
                        fftRB <= data_in;
                        addr <= idxBaixo + 1024;
                        state <= WAIT_DATA4;
                    end
                WAIT_DATA4:
                    state <= READ_MEM4;
                READ_MEM4:
                    begin
                        fftIB <= data_in;
                        state <= MULT1;
                    end
                MULT1:
                    begin
                        if(LOOP_1_Counter == 3 && LOOP_2_Counter == 1 && LOOP_3_Counter == 2) begin
                            $display("fftRB: %d WnI: %d fftIB: %d WnR: %d", fftRB, WnI_op, fftIB, WnR_op);
                        end
                        temp2R_aux <= ((fftRB * WnR_op) - (fftIB * WnI_op));
                        temp2I_aux <= ((fftRB * WnI_op) + (fftIB * WnR_op));
                        state <= MULT2;
                    end
                MULT2:
                    begin
                        fftRB <= temp2R;
                        fftIB <= temp2I;
                        state <= MULT3;
                    end
                MULT3:
                    begin
                        fftRC <= fftRC + fftRB;
                        fftIC <= fftIC + fftIB;
                        state <= MULT4;
                    end
                MULT4:
                    begin
                        fftRB <= fftRB - tempR;
                        fftIB <= fftIB - tempI;
                        state <= DIV;
                    end
                DIV:
                    begin
                        fftRC <= fftRC / 2;
                        fftIC <= fftIC / 2;
                        fftRB <= fftRB / 2;
                        fftIB <= fftIB / 2;
                        state <= STORE1;
                    end
                STORE1:
                    begin
                        // if(LOOP_1_Counter == 2) begin
                        //     $display("%d \t fftRC: %d fftIC: %d fftRB: %d fftIB: %d",debug_count, fftRC, fftIC, fftRB, fftIB);
                        //     debug_count = debug_count + 1;
                        // end
                        write_enable <= 1;
                        addr <= idxCima;
                        data_out <= fftRC;
                        state <= STORE2;
                    end
                STORE2:
                    begin
                        addr <= idxCima + 1024;
                        data_out <= fftIC;
                        state <= STORE3;
                    end
                STORE3:
                    begin
                        addr <= idxBaixo;
                        data_out <= fftRB;
                        state <= STORE4;
                    end
                STORE4:
                    begin
                        addr <= idxBaixo + 1024;
                        data_out <= fftIB;
                        state <= LOOP_3;
                    end
                END:
                    begin
                        state <= END;                        
                        fft_done <= 1;
                    end
                default:
                    state <= IDLE;
            endcase
        end
    end

endmodule